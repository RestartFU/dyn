module rsh

